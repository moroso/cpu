parameter EXN_CODE_NOERR = 5'b0;
parameter EXN_CODE_INST_PF = 5'b00001;
parameter EXN_CODE_ILL = 5'b00010;
parameter EXN_CODE_NO_PERM = 5'b00011;
parameter EXN_CODE_DUP_DEST = 5'b00100;
parameter EXN_CODE_DATA_PF = 5'b00101;
parameter EXN_CODE_BAD_PHYSADDR = 5'b00110;
parameter EXN_CODE_DIVZERO = 5'b00111;
parameter EXN_CODE_INTERRUPT = 5'b01000;
parameter EXN_CODE_SYSCALL = 5'b01001;
parameter EXN_CODE_BREAK = 5'b01010;
