parameter OPER_TYPE_ALU = 2'b000;
parameter OPER_TYPE_BRANCH = 2'b001;
parameter OPER_TYPE_LSU = 2'b010;
parameter OPER_TYPE_OTHER = 2'b11;
