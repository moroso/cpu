
parameter OPCODE_ERET = 9'b