parameter OPER_TYPE_ALU = 2'b00;
parameter OPER_TYPE_BRANCH = 2'b01;
parameter OPER_TYPE_LSU = 2'b10;
parameter OPER_TYPE_OTHER = 2'b11;
