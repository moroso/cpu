parameter LTC_OPC_READ         = 3'b000;
parameter LTC_OPC_WRITE        = 3'b001;
parameter LTC_OPC_READTHROUGH  = 3'b010;
parameter LTC_OPC_WRITETHROUGH = 3'b011;
parameter LTC_OPC_PREFETCH     = 3'b100;
parameter LTC_OPC_CLEAN        = 3'b110;
