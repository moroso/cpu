// Flag bit offsets for page tables.
parameter PAGETAB_PRESENT = 0;
parameter PAGETAB_WRITEABLE = 1;
parameter PAGETAB_KERNEL = 2;
parameter PAGETAB_GLOBAL = 3;
