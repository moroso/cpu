parameter COPROC_OP_BREAK = 4'b0001;
parameter COPROC_OP_SYSCALL = 4'b0010;
parameter COPROC_OP_FENCE = 4'b0011;
parameter COPROC_OP_ERET = 4'b0100;
parameter COPROC_OP_FLUSH = 4'b0101;
parameter COPROC_OP_MFC = 4'b0110;
parameter COPROC_OP_MTC = 4'b0111;
parameter COPROC_OP_MULT = 4'b1000;
parameter COPROC_OP_DIV = 4'b1001;
parameter COPROC_OP_MFHI = 4'b1010;
parameter COPROC_OP_MTHI = 4'b1011;
